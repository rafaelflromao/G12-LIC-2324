    Mac OS X            	   2   �      �                                      ATTR       �   �   H                  �   H  com.apple.macl    �}Z�Y
J���N/��p                                                      