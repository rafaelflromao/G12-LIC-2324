    Mac OS X            	   2   �                                           ATTR         �   X                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl   MXf    �w�
     �}Z�Y
J���N/��p                                                      