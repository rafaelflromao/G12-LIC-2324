    Mac OS X            	   2  �     �                                      ATTR      �   �   �                  �   �  "com.apple.LaunchServices.OpenWith      ~     com.apple.lastuseddate#PS      �   H  com.apple.macl   bplist00�WversionTpath_bundleidentifier _ /Applications/DevOp/Brackets.app_io.brackets.appshell/1T                            kzVf    �!     �}Z�Y
J���N/��p                                                      